module top (
  input  logic clk
);
  // TODO: your design here
endmodule
